module XOR2(A, B, Cout);
  input A, B;
  output Cout;
  
  assign Cout = A ^ B; // Cout = A XOR B
  
endmodule